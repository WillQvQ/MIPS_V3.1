`timescale 1ns / 1ps

module hazardunit(
    
);
    
endmodule